--
-- Pixel generation circuit
-- (c) OptimalBits Sweden AB 2015.
--


